library IEEE;
use IEEE.std_logic_1164.all;

entity GeradorTick is
	port (
		clock						: in  std_logic;
		reset						: in  std_logic;
		tick						: out std_logic
	);
end GeradorTick;

architecture hierarquica of GeradorTick is





begin



end hierarquica;
