library IEEE;
use IEEE.std_logic_1164.all;

entity fluxo_dados is
  port ();
end fluxo_dados;

architecture combinatorio of fluxo_dados is

begin


end combinatorio;
