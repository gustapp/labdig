library IEEE;
use IEEE.std_logic_1164.all;

entity RecepcaoSerial is
  port (
    clock     : in std_logic;
    dados     : out std_logic
  );
end RecepcaoSerial;

architecture hierarquico of RecepcaoSerial is

begin


end hierarquico;
